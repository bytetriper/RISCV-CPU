`include "Icache.v"
module TEST();
    
endmodule