module Fetcher();
endmodule
