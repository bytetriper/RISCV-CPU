module ICache();
endmodule
